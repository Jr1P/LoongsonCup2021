`timescale 1ns/1ps

// * Pipeline stall and refresh
module cu(
    input   
    input


    output  if_id_stall,
    output  id_ex_stall,
    output  ex_mem_stall,
    output  mem_wb_stall,

    output  if_id_refresh,
    output  id_ex_refresh,
    output  ex_mem_refresh,
    output  mem_wb_refresh
);



endmodule
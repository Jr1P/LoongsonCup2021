`timescale 1ns/1ps

module pc(

);

always @(posedge clk) begin

end

endmodule
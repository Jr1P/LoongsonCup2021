`timescale 1ns/1ps

module pc(

);
// TODO:
always @(posedge clk) begin

end

endmodule
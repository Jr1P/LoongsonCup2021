`timescale 1ns/1ps

module cu(

    output 
);



endmodule
`timescale 1ns/1ps

module cu(

);

always @(posedge clk) begin

end

endmodule